LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

ENTITY decod7seg IS
	PORT (
		c : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		h : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END decod7seg;
ARCHITECTURE decoder OF decod7seg IS
BEGIN
	h <=  "1000000" WHEN c = "0000" ELSE --0
	"1111001" WHEN c = "0001" ELSE --1
	"0100100" WHEN c = "0010" ELSE --2
	"0110000" WHEN c = "0011" ELSE --3
	"0011001" WHEN c = "0100" ELSE --4
	"0010010" WHEN c = "0101" ELSE --5
	"0000010" WHEN c = "0110" ELSE --6
	"1111000" WHEN c = "0111" ELSE --7
	"0000000" WHEN c = "1000" ELSE --8
	"0010000" WHEN c = "1001" ELSE --9
	"0001000" WHEN c = "1010" ELSE --A
	"0000011" WHEN c = "1011" ELSE --b
	"1000110" WHEN c = "1100" ELSE --c
	"0100001" WHEN c = "1101" ELSE --d
	"0000110" WHEN c = "1110" ELSE --E
	"0001110"; --F
END decoder;